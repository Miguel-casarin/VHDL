library ieee;
use ieee.std_logic_1164.all;

entity r_or is
    port(
        a, b : in std_logic;
        y : out std_logic);
end r_or;

architecture c_or of r_or is

begin
    y <= a or b;
end c_or; 